7890
htns
1234
